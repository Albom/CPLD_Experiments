module Button (button, LED, clk);

input button;
output LED;
input clk;

initial begin

end


assign LED = button;

endmodule 